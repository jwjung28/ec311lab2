module display_control ();

endmodule
