module clock_divider ();

endmodule
