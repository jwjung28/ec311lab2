module top (
    input clock, reset, mode_select, increment,
    output [3:0] digit_select,
    output [6:0] seg
    );

endmodule
