module counter_8bit (
    input clock, reset, increment,
    output [7:0] count
    );

endmodule