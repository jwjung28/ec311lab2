module counter16 ();

endmodule
