module seven_seg_decoder ();

endmodule
